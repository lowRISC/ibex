// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

class dv_base_virtual_sequencer #(
  type CFG_T = dv_base_env_cfg,
  type COV_T = dv_base_env_cov
) extends uvm_sequencer;
  `uvm_component_param_utils(dv_base_virtual_sequencer#(CFG_T, COV_T))

  CFG_T cfg;
  COV_T cov;

  `uvm_component_new

endclass
