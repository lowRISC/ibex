// Copyright lowRISC contributors (OpenTitan project).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//

package rv_dm_pkg;

  parameter int NrHarts = 1;

  typedef logic [31:0] next_dm_addr_t;

  parameter next_dm_addr_t NEXT_DM_ADDR_DEFAULT = '0;

endpackage : rv_dm_pkg
