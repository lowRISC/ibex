// Copyleft ISOLDE 2025

package isolde_soc_package;

  parameter int unsigned DEFAULT_DW = 32; // Default Data Width
  parameter int unsigned DEFAULT_AW = 32; // Default Address Width
  parameter int unsigned DEFAULT_BW = 8;  // Default Byte Width
  parameter int unsigned DEFAULT_WW = 32; // Default Word Width
  parameter int unsigned DEFAULT_UW = 0;  // Default User Width



endpackage // isolde_soc_package
