// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//

package top_pkg;

localparam int TL_AW=32;
localparam int TL_DW=32;    // = TL_DBW * 8; TL_DBW must be a power-of-two
localparam int TL_AIW=8;    // a_source, d_source
localparam int TL_DIW=1;    // d_sink
localparam int TL_DUW=16;   // d_user
localparam int TL_DBW=(TL_DW>>3);
localparam int TL_SZW=$clog2($clog2(TL_DBW)+1);
localparam int FLASH_BANKS=2;
localparam int FLASH_PAGES_PER_BANK=256;
localparam int FLASH_WORDS_PER_PAGE=256;
localparam int FLASH_BYTES_PER_WORD=4;
localparam int FLASH_BKW = $clog2(FLASH_BANKS);
localparam int FLASH_PGW = $clog2(FLASH_PAGES_PER_BANK);
localparam int FLASH_WDW = $clog2(FLASH_WORDS_PER_PAGE);
localparam int FLASH_AW = FLASH_BKW + FLASH_PGW + FLASH_WDW;
localparam int FLASH_DW = FLASH_BYTES_PER_WORD * 8;

endpackage
